VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM32
  CLASS BLOCK ;
  FOREIGN RAM32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 401.580 BY 136.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 17.720 401.580 18.320 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 29.960 401.580 30.560 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 42.200 401.580 42.800 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 54.440 401.580 55.040 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 66.680 401.580 67.280 ;
    END
  END A0[4]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 399.580 78.920 401.580 79.520 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 7.910 134.000 8.190 136.000 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 134.000 132.390 136.000 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 134.000 144.810 136.000 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 156.950 134.000 157.230 136.000 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 169.370 134.000 169.650 136.000 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 134.000 182.070 136.000 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 194.210 134.000 194.490 136.000 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 206.630 134.000 206.910 136.000 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 134.000 219.330 136.000 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 231.470 134.000 231.750 136.000 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 243.890 134.000 244.170 136.000 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 20.330 134.000 20.610 136.000 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 256.310 134.000 256.590 136.000 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 268.730 134.000 269.010 136.000 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 281.150 134.000 281.430 136.000 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 293.570 134.000 293.850 136.000 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 305.990 134.000 306.270 136.000 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 318.410 134.000 318.690 136.000 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 330.830 134.000 331.110 136.000 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 343.250 134.000 343.530 136.000 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 355.670 134.000 355.950 136.000 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 368.090 134.000 368.370 136.000 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 32.750 134.000 33.030 136.000 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 380.510 134.000 380.790 136.000 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 134.000 393.210 136.000 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 134.000 45.450 136.000 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 57.590 134.000 57.870 136.000 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 70.010 134.000 70.290 136.000 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 82.430 134.000 82.710 136.000 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 134.000 95.130 136.000 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 107.270 134.000 107.550 136.000 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 134.000 119.970 136.000 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 5.480 401.580 6.080 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 133.520 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 133.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 133.520 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 91.160 401.580 91.760 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 103.400 401.580 104.000 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 115.640 401.580 116.240 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 399.580 127.880 401.580 128.480 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 2.570 129.145 399.010 131.975 ;
        RECT 2.570 123.705 399.010 126.535 ;
        RECT 2.570 118.265 399.010 121.095 ;
        RECT 2.570 112.825 399.010 115.655 ;
        RECT 2.570 107.435 399.010 110.215 ;
        RECT 2.570 107.385 84.715 107.435 ;
        RECT 2.570 104.725 85.175 104.775 ;
        RECT 2.570 101.995 399.010 104.725 ;
        RECT 2.570 101.945 84.715 101.995 ;
        RECT 2.570 99.285 85.175 99.335 ;
        RECT 2.570 96.555 399.010 99.285 ;
        RECT 2.570 96.505 84.715 96.555 ;
        RECT 2.570 93.845 85.175 93.895 ;
        RECT 2.570 91.115 399.010 93.845 ;
        RECT 2.570 91.065 84.715 91.115 ;
        RECT 2.570 88.405 85.175 88.455 ;
        RECT 2.570 85.675 399.010 88.405 ;
        RECT 2.570 85.625 84.715 85.675 ;
        RECT 2.570 82.965 85.175 83.015 ;
        RECT 2.570 80.235 399.010 82.965 ;
        RECT 2.570 80.185 84.715 80.235 ;
        RECT 2.570 77.525 85.175 77.575 ;
        RECT 2.570 74.795 399.010 77.525 ;
        RECT 2.570 74.745 84.715 74.795 ;
        RECT 2.570 72.085 85.175 72.135 ;
        RECT 2.570 69.355 399.010 72.085 ;
        RECT 2.570 69.305 84.715 69.355 ;
        RECT 2.570 66.645 85.175 66.695 ;
        RECT 2.570 63.865 399.010 66.645 ;
        RECT 2.570 58.425 399.010 61.255 ;
        RECT 2.570 52.985 399.010 55.815 ;
        RECT 2.570 47.595 399.010 50.375 ;
        RECT 2.570 47.545 84.715 47.595 ;
        RECT 2.570 44.885 85.175 44.935 ;
        RECT 2.570 42.155 399.010 44.885 ;
        RECT 2.570 42.105 84.715 42.155 ;
        RECT 2.570 39.445 85.175 39.495 ;
        RECT 2.570 36.715 399.010 39.445 ;
        RECT 2.570 36.665 84.715 36.715 ;
        RECT 2.570 34.005 85.175 34.055 ;
        RECT 2.570 31.275 399.010 34.005 ;
        RECT 2.570 31.225 84.715 31.275 ;
        RECT 2.570 28.565 85.175 28.615 ;
        RECT 2.570 25.835 399.010 28.565 ;
        RECT 2.570 25.785 84.715 25.835 ;
        RECT 2.570 23.125 85.175 23.175 ;
        RECT 2.570 20.395 399.010 23.125 ;
        RECT 2.570 20.345 84.715 20.395 ;
        RECT 2.570 17.685 85.175 17.735 ;
        RECT 2.570 14.955 399.010 17.685 ;
        RECT 2.570 14.905 84.715 14.955 ;
        RECT 2.570 12.245 85.175 12.295 ;
        RECT 2.570 9.515 399.010 12.245 ;
        RECT 2.570 9.465 84.715 9.515 ;
        RECT 2.570 6.805 85.175 6.855 ;
        RECT 2.570 4.025 399.010 6.805 ;
      LAYER li1 ;
        RECT 2.760 2.635 398.820 133.365 ;
      LAYER met1 ;
        RECT 2.760 0.040 398.820 135.960 ;
      LAYER met2 ;
        RECT 3.310 133.720 7.630 135.990 ;
        RECT 8.470 133.720 20.050 135.990 ;
        RECT 20.890 133.720 32.470 135.990 ;
        RECT 33.310 133.720 44.890 135.990 ;
        RECT 45.730 133.720 57.310 135.990 ;
        RECT 58.150 133.720 69.730 135.990 ;
        RECT 70.570 133.720 82.150 135.990 ;
        RECT 82.990 133.720 94.570 135.990 ;
        RECT 95.410 133.720 106.990 135.990 ;
        RECT 107.830 133.720 119.410 135.990 ;
        RECT 120.250 133.720 131.830 135.990 ;
        RECT 132.670 133.720 144.250 135.990 ;
        RECT 145.090 133.720 156.670 135.990 ;
        RECT 157.510 133.720 169.090 135.990 ;
        RECT 169.930 133.720 181.510 135.990 ;
        RECT 182.350 133.720 193.930 135.990 ;
        RECT 194.770 133.720 206.350 135.990 ;
        RECT 207.190 133.720 218.770 135.990 ;
        RECT 219.610 133.720 231.190 135.990 ;
        RECT 232.030 133.720 243.610 135.990 ;
        RECT 244.450 133.720 256.030 135.990 ;
        RECT 256.870 133.720 268.450 135.990 ;
        RECT 269.290 133.720 280.870 135.990 ;
        RECT 281.710 133.720 293.290 135.990 ;
        RECT 294.130 133.720 305.710 135.990 ;
        RECT 306.550 133.720 318.130 135.990 ;
        RECT 318.970 133.720 330.550 135.990 ;
        RECT 331.390 133.720 342.970 135.990 ;
        RECT 343.810 133.720 355.390 135.990 ;
        RECT 356.230 133.720 367.810 135.990 ;
        RECT 368.650 133.720 380.230 135.990 ;
        RECT 381.070 133.720 392.650 135.990 ;
        RECT 393.490 133.720 398.270 135.990 ;
        RECT 3.310 2.280 398.270 133.720 ;
        RECT 3.310 0.010 7.630 2.280 ;
        RECT 8.470 0.010 20.050 2.280 ;
        RECT 20.890 0.010 32.470 2.280 ;
        RECT 33.310 0.010 44.890 2.280 ;
        RECT 45.730 0.010 57.310 2.280 ;
        RECT 58.150 0.010 69.730 2.280 ;
        RECT 70.570 0.010 82.150 2.280 ;
        RECT 82.990 0.010 94.570 2.280 ;
        RECT 95.410 0.010 106.990 2.280 ;
        RECT 107.830 0.010 119.410 2.280 ;
        RECT 120.250 0.010 131.830 2.280 ;
        RECT 132.670 0.010 144.250 2.280 ;
        RECT 145.090 0.010 156.670 2.280 ;
        RECT 157.510 0.010 169.090 2.280 ;
        RECT 169.930 0.010 181.510 2.280 ;
        RECT 182.350 0.010 193.930 2.280 ;
        RECT 194.770 0.010 206.350 2.280 ;
        RECT 207.190 0.010 218.770 2.280 ;
        RECT 219.610 0.010 231.190 2.280 ;
        RECT 232.030 0.010 243.610 2.280 ;
        RECT 244.450 0.010 256.030 2.280 ;
        RECT 256.870 0.010 268.450 2.280 ;
        RECT 269.290 0.010 280.870 2.280 ;
        RECT 281.710 0.010 293.290 2.280 ;
        RECT 294.130 0.010 305.710 2.280 ;
        RECT 306.550 0.010 318.130 2.280 ;
        RECT 318.970 0.010 330.550 2.280 ;
        RECT 331.390 0.010 342.970 2.280 ;
        RECT 343.810 0.010 355.390 2.280 ;
        RECT 356.230 0.010 367.810 2.280 ;
        RECT 368.650 0.010 380.230 2.280 ;
        RECT 381.070 0.010 392.650 2.280 ;
        RECT 393.490 0.010 398.270 2.280 ;
      LAYER met3 ;
        RECT 3.285 128.880 399.580 135.825 ;
        RECT 3.285 127.480 399.180 128.880 ;
        RECT 3.285 116.640 399.580 127.480 ;
        RECT 3.285 115.240 399.180 116.640 ;
        RECT 3.285 104.400 399.580 115.240 ;
        RECT 3.285 103.000 399.180 104.400 ;
        RECT 3.285 92.160 399.580 103.000 ;
        RECT 3.285 90.760 399.180 92.160 ;
        RECT 3.285 79.920 399.580 90.760 ;
        RECT 3.285 78.520 399.180 79.920 ;
        RECT 3.285 67.680 399.580 78.520 ;
        RECT 3.285 66.280 399.180 67.680 ;
        RECT 3.285 55.440 399.580 66.280 ;
        RECT 3.285 54.040 399.180 55.440 ;
        RECT 3.285 43.200 399.580 54.040 ;
        RECT 3.285 41.800 399.180 43.200 ;
        RECT 3.285 30.960 399.580 41.800 ;
        RECT 3.285 29.560 399.180 30.960 ;
        RECT 3.285 18.720 399.580 29.560 ;
        RECT 3.285 17.320 399.180 18.720 ;
        RECT 3.285 6.480 399.580 17.320 ;
        RECT 3.285 5.080 399.180 6.480 ;
        RECT 3.285 0.175 399.580 5.080 ;
      LAYER met4 ;
        RECT 164.975 17.855 171.480 112.025 ;
        RECT 173.880 17.855 248.280 112.025 ;
        RECT 250.680 17.855 325.080 112.025 ;
        RECT 327.480 17.855 391.625 112.025 ;
  END
END RAM32
END LIBRARY

